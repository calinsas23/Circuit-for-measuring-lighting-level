** Profile: "SCHEMATIC1-monte"  [ D:\Homeworks\An 2 sem 2\Tehnici CAD\Proiect-final\Final-Corect\proiect_cad-PSpiceFiles\SCHEMATIC1\monte.sim ] 

** Creating circuit file "monte.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of D:\Homeworks\An 2 sem 2\Tehnici CAD\Projects\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "D:\Homeworks\An 2 sem 2\Tehnici CAD\Proiect-final\Final-Corect\leduri.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.WCASE TRAN v([LED]) YMAX VARY BOTH  HI 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
