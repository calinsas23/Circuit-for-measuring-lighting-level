** Profile: "SCHEMATIC1-dc"  [ D:\Homeworks\An 2 sem 2\Tehnici CAD\Proiect-final\Final-Corect\proiect_cad-pspicefiles\schematic1\dc.sim ] 

** Creating circuit file "dc.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of D:\Homeworks\An 2 sem 2\Tehnici CAD\Projects\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "D:\Homeworks\An 2 sem 2\Tehnici CAD\Proiect-final\Final-Corect\leduri.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.MC 10 TRAN v([LED]) YMAX OUTPUT ALL SEED=200 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
